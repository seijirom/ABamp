* Created by KLayout

* cell amp_ab
.SUBCKT amp_ab
* net 28 SUBSTRATE
* device instance $1 m0 *1 213.34,-155.03 NMOS
M$1 4 1 28 28 NMOS L=1U W=8000U AS=8160P AD=8160P PS=8364U PD=8364U
* device instance $101 r0 *1 146.39,15.36 PMOS
M$101 3 6 7 3 PMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $105 r0 *1 134.39,-31.64 NMOS
M$105 1 14 7 28 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $106 m90 *1 124.39,-31.64 NMOS
M$106 9 14 14 28 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $107 m90 *1 88.89,-32.14 CAP
C$107 10 7 1.04e-11 CAP
* device instance $108 m90 *1 148.39,-31.64 PMOS
M$108 7 11 1 7 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $109 r0 *1 164.39,-31.64 PMOS
M$109 15 11 11 15 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $110 r0 *1 20.39,2.86 HRES
R$110 5 3 120750 HRES
* device instance $111 r0 *1 -1.11,-34.64 HRES
R$111 3 8 20000 HRES
* device instance $112 r0 *1 9.39,-34.64 HRES
R$112 28 8 20000 HRES
* device instance $113 m90 *1 52.39,-44.14 NMOS
M$113 12 2 10 28 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $114 r180 *1 52.39,-23.14 NMOS
M$114 6 2 10 28 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $115 r0 *1 34.39,-44.14 NMOS
M$115 12 8 13 28 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $116 m0 *1 34.39,-23.14 NMOS
M$116 17 8 13 28 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $117 m0 *1 127.39,-78.64 NMOS
M$117 1 5 28 28 NMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $121 m0 *1 34.39,-78.64 NMOS
M$121 12 5 28 28 NMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $125 r180 *1 1.39,-78.64 NMOS
M$125 16 5 28 28 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $127 r180 *1 21.39,-78.64 NMOS
M$127 5 5 28 28 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $129 m0 *1 160.89,-79.14 NMOS
M$129 11 5 28 28 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $131 r0 *1 -3.61,14.86 PMOS
M$131 3 16 16 3 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $133 m90 *1 58.89,14.86 PMOS
M$133 3 17 6 3 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $135 r0 *1 122.89,15.36 PMOS
M$135 3 16 14 3 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $137 r0 *1 34.89,14.86 PMOS
M$137 3 17 17 3 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $140 m90 *1 141.91,117.55 HRES
R$140 29 2 10000 HRES
* device instance $148 m90 *1 191.91,147.55 HRES
R$148 4 2 110000 HRES
* device instance $151 r0 *1 214.49,-28.01 PMOS
M$151 3 7 4 3 PMOS L=1U W=28000U AS=28560P AD=28560P PS=28968U PD=28968U
* device instance $351 r180 *1 78.67,85.35 PMOS
M$351 3 15 15 3 PMOS L=1U W=1280U AS=1320P AD=1320P PS=1386U PD=1386U
* device instance $383 m90 *1 77.02,138.26 NMOS
M$383 28 9 9 28 NMOS L=1U W=1280U AS=1320P AD=1320P PS=1386U PD=1386U
.ENDS amp_ab
