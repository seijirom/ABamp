* Created by KLayout

* cell amp_ab
.SUBCKT amp_ab
* net 28 SUBSTRATE
* cell instance $2 m90 *1 56.39,-51.14
X$2 11 9 1 28 Nch$5
* cell instance $3 r180 *1 56.39,-16.14
X$3 5 9 1 28 Nch$5
* cell instance $7 r0 *1 211.99,-101.01
X$7 3 6 2 2 Pch$6
* cell instance $8 r0 *1 371.99,-101.01
X$8 3 6 2 2 Pch$6
* cell instance $9 r180 *1 81.17,108.35
X$9 2 2 2 2 Pch$7
* cell instance $10 r0 *1 -7.61,-8.14
X$10 2 15 15 2 Pch$2
* cell instance $11 r0 *1 142.39,-7.64
X$11 6 5 2 2 Pch$4
* cell instance $12 m90 *1 62.89,-8.14
X$12 2 5 16 2 Pch$2
* cell instance $13 r0 *1 118.89,-7.64
X$13 2 14 15 2 Pch$2
* cell instance $14 r0 *1 30.89,-8.14
X$14 2 16 16 2 Pch$2
* cell instance $15 r0 *1 160.39,-44.64
X$15 2 10 10 2 Pch$5
* cell instance $16 r180 *1 523.93,195.89
X$16 2 6 3 2 Pch$6
* cell instance $17 r180 *1 363.75,195.99
X$17 2 6 3 2 Pch$6
* cell instance $22 m90 *1 112.89,-82.14
X$22 6 9 Capacitor$1
* cell instance $23 m0 *1 210.84,-112.03
X$23 3 28 28 28 Nch$7
* cell instance $24 m0 *1 372.95,-112.05
X$24 3 28 28 28 Nch$7
* cell instance $26 m0 *1 30.39,-55.64
X$26 11 28 4 28 Nch$3
* cell instance $27 r180 *1 5.39,-55.64
X$27 15 28 4 28 Nch$1
* cell instance $28 r180 *1 25.39,-55.64
X$28 4 28 4 28 Nch$1
* cell instance $29 m0 *1 123.39,-55.64
X$29 13 28 4 28 Nch$3
* cell instance $30 m0 *1 156.89,-56.14
X$30 10 28 4 28 Nch$1
* cell instance $31 m90 *1 152.39,-44.64
X$31 6 28 10 6 Pch$5
* cell instance $32 r0 *1 130.39,-44.64
X$32 13 6 14 28 Nch$4
* cell instance $37 r0 *1 30.39,-51.14
X$37 11 12 7 28 Nch$5
* cell instance $38 m0 *1 30.39,-16.14
X$38 16 12 7 28 Nch$5
* cell instance $40 m90 *1 128.39,-44.64
X$40 8 14 14 28 Nch$4
* cell instance $41 m90 *1 79.52,115.26
X$41 28 8 8 28 Nch$6
* device instance $1 r0 *1 -1.11,-34.64 HRES
R$1 2 7 20000
* device instance $2 r0 *1 9.39,-34.64 HRES
R$2 28 7 20000
* device instance $3 r0 *1 20.39,2.86 HRES
R$3 4 2 120750
* device instance $4 r0 *1 116.91,87.55 HRES
R$4 17 21 10000
* device instance $5 r0 *1 141.91,87.55 HRES
R$5 18 17 10000
* device instance $6 r0 *1 166.91,87.55 HRES
R$6 18 20 10000
* device instance $7 r0 *1 191.91,87.55 HRES
R$7 3 19 10000
* device instance $8 r0 *1 116.91,117.55 HRES
R$8 21 23 10000
* device instance $9 r0 *1 141.91,117.55 HRES
R$9 1 25 10000
* device instance $10 r0 *1 166.91,117.55 HRES
R$10 20 26 10000
* device instance $11 r0 *1 191.91,117.55 HRES
R$11 19 22 10000
* device instance $12 r0 *1 116.91,147.55 HRES
R$12 23 24 10000
* device instance $13 r0 *1 141.91,147.55 HRES
R$13 25 24 10000
* device instance $14 r0 *1 166.91,147.55 HRES
R$14 26 27 10000
* device instance $15 r0 *1 191.91,147.55 HRES
R$15 22 27 10000
.ENDS amp_ab

* cell Pch$4
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch$4 1 2 3 4
* device instance $1 r0 *1 4,23 PMOS
M$1 3 2 1 4 PMOS L=4U W=40U AS=80P AD=40P PS=84U PD=42U
* device instance $2 r0 *1 10,23 PMOS
M$2 1 2 3 4 PMOS L=4U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $3 r0 *1 16,23 PMOS
M$3 3 2 1 4 PMOS L=4U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $4 r0 *1 22,23 PMOS
M$4 1 2 3 4 PMOS L=4U W=40U AS=40P AD=80P PS=42U PD=84U
.ENDS Pch$4

* cell Nch$4
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$4 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 4,13 NMOS
M$1 1 3 2 4 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS Nch$4

* cell Nch$7
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$7 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 2.5,23 NMOS
M$1 1 3 2 4 NMOS L=1U W=40U AS=80P AD=40P PS=84U PD=42U
* device instance $2 r0 *1 5.5,23 NMOS
M$2 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $3 r0 *1 8.5,23 NMOS
M$3 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $4 r0 *1 11.5,23 NMOS
M$4 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $5 r0 *1 14.5,23 NMOS
M$5 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $6 r0 *1 17.5,23 NMOS
M$6 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $7 r0 *1 20.5,23 NMOS
M$7 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $8 r0 *1 23.5,23 NMOS
M$8 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $9 r0 *1 26.5,23 NMOS
M$9 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $10 r0 *1 29.5,23 NMOS
M$10 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $11 r0 *1 32.5,23 NMOS
M$11 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $12 r0 *1 35.5,23 NMOS
M$12 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $13 r0 *1 38.5,23 NMOS
M$13 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $14 r0 *1 41.5,23 NMOS
M$14 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $15 r0 *1 44.5,23 NMOS
M$15 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $16 r0 *1 47.5,23 NMOS
M$16 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $17 r0 *1 50.5,23 NMOS
M$17 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $18 r0 *1 53.5,23 NMOS
M$18 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $19 r0 *1 56.5,23 NMOS
M$19 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $20 r0 *1 59.5,23 NMOS
M$20 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $21 r0 *1 62.5,23 NMOS
M$21 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $22 r0 *1 65.5,23 NMOS
M$22 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $23 r0 *1 68.5,23 NMOS
M$23 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $24 r0 *1 71.5,23 NMOS
M$24 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $25 r0 *1 74.5,23 NMOS
M$25 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $26 r0 *1 77.5,23 NMOS
M$26 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $27 r0 *1 80.5,23 NMOS
M$27 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $28 r0 *1 83.5,23 NMOS
M$28 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $29 r0 *1 86.5,23 NMOS
M$29 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $30 r0 *1 89.5,23 NMOS
M$30 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $31 r0 *1 92.5,23 NMOS
M$31 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $32 r0 *1 95.5,23 NMOS
M$32 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $33 r0 *1 98.5,23 NMOS
M$33 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $34 r0 *1 101.5,23 NMOS
M$34 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $35 r0 *1 104.5,23 NMOS
M$35 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $36 r0 *1 107.5,23 NMOS
M$36 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $37 r0 *1 110.5,23 NMOS
M$37 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $38 r0 *1 113.5,23 NMOS
M$38 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $39 r0 *1 116.5,23 NMOS
M$39 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $40 r0 *1 119.5,23 NMOS
M$40 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $41 r0 *1 122.5,23 NMOS
M$41 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $42 r0 *1 125.5,23 NMOS
M$42 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $43 r0 *1 128.5,23 NMOS
M$43 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $44 r0 *1 131.5,23 NMOS
M$44 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $45 r0 *1 134.5,23 NMOS
M$45 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $46 r0 *1 137.5,23 NMOS
M$46 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $47 r0 *1 140.5,23 NMOS
M$47 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $48 r0 *1 143.5,23 NMOS
M$48 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $49 r0 *1 146.5,23 NMOS
M$49 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $50 r0 *1 149.5,23 NMOS
M$50 2 3 1 4 NMOS L=1U W=40U AS=40P AD=80P PS=42U PD=84U
.ENDS Nch$7

* cell Capacitor$1
* pin 
* pin 
.SUBCKT Capacitor$1 1 2
* device instance $1 r0 *1 24,50 CAP
C$1 2 1 1.04e-11
.ENDS Capacitor$1

* cell Pch$5
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch$5 1 2 3 4
* device instance $1 r0 *1 4,13 PMOS
M$1 1 3 2 4 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS Pch$5

* cell Nch$5
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$5 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 4,7 NMOS
M$1 1 3 2 4 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
.ENDS Nch$5

* cell Nch$3
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$3 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 4,23 NMOS
M$1 1 3 2 4 NMOS L=4U W=40U AS=80P AD=40P PS=84U PD=42U
* device instance $2 r0 *1 10,23 NMOS
M$2 2 3 1 4 NMOS L=4U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $3 r0 *1 16,23 NMOS
M$3 1 3 2 4 NMOS L=4U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $4 r0 *1 22,23 NMOS
M$4 2 3 1 4 NMOS L=4U W=40U AS=40P AD=80P PS=42U PD=84U
.ENDS Nch$3

* cell Nch$1
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$1 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 4,23 NMOS
M$1 1 3 2 4 NMOS L=4U W=40U AS=80P AD=40P PS=84U PD=42U
* device instance $2 r0 *1 10,23 NMOS
M$2 2 3 1 4 NMOS L=4U W=40U AS=40P AD=80P PS=42U PD=84U
.ENDS Nch$1

* cell Pch$2
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch$2 1 2 3 4
* device instance $1 r0 *1 4,23 PMOS
M$1 1 3 2 4 PMOS L=4U W=40U AS=80P AD=40P PS=84U PD=42U
* device instance $2 r0 *1 10,23 PMOS
M$2 2 3 1 4 PMOS L=4U W=40U AS=40P AD=80P PS=42U PD=84U
.ENDS Pch$2

* cell Pch$6
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch$6 1 2 3 4
* device instance $1 r0 *1 2.5,73 PMOS
M$1 3 2 1 4 PMOS L=1U W=140U AS=280P AD=140P PS=284U PD=142U
* device instance $2 r0 *1 5.5,73 PMOS
M$2 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $3 r0 *1 8.5,73 PMOS
M$3 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $4 r0 *1 11.5,73 PMOS
M$4 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $5 r0 *1 14.5,73 PMOS
M$5 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $6 r0 *1 17.5,73 PMOS
M$6 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $7 r0 *1 20.5,73 PMOS
M$7 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $8 r0 *1 23.5,73 PMOS
M$8 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $9 r0 *1 26.5,73 PMOS
M$9 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $10 r0 *1 29.5,73 PMOS
M$10 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $11 r0 *1 32.5,73 PMOS
M$11 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $12 r0 *1 35.5,73 PMOS
M$12 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $13 r0 *1 38.5,73 PMOS
M$13 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $14 r0 *1 41.5,73 PMOS
M$14 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $15 r0 *1 44.5,73 PMOS
M$15 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $16 r0 *1 47.5,73 PMOS
M$16 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $17 r0 *1 50.5,73 PMOS
M$17 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $18 r0 *1 53.5,73 PMOS
M$18 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $19 r0 *1 56.5,73 PMOS
M$19 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $20 r0 *1 59.5,73 PMOS
M$20 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $21 r0 *1 62.5,73 PMOS
M$21 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $22 r0 *1 65.5,73 PMOS
M$22 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $23 r0 *1 68.5,73 PMOS
M$23 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $24 r0 *1 71.5,73 PMOS
M$24 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $25 r0 *1 74.5,73 PMOS
M$25 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $26 r0 *1 77.5,73 PMOS
M$26 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $27 r0 *1 80.5,73 PMOS
M$27 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $28 r0 *1 83.5,73 PMOS
M$28 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $29 r0 *1 86.5,73 PMOS
M$29 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $30 r0 *1 89.5,73 PMOS
M$30 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $31 r0 *1 92.5,73 PMOS
M$31 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $32 r0 *1 95.5,73 PMOS
M$32 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $33 r0 *1 98.5,73 PMOS
M$33 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $34 r0 *1 101.5,73 PMOS
M$34 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $35 r0 *1 104.5,73 PMOS
M$35 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $36 r0 *1 107.5,73 PMOS
M$36 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $37 r0 *1 110.5,73 PMOS
M$37 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $38 r0 *1 113.5,73 PMOS
M$38 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $39 r0 *1 116.5,73 PMOS
M$39 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $40 r0 *1 119.5,73 PMOS
M$40 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $41 r0 *1 122.5,73 PMOS
M$41 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $42 r0 *1 125.5,73 PMOS
M$42 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $43 r0 *1 128.5,73 PMOS
M$43 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $44 r0 *1 131.5,73 PMOS
M$44 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $45 r0 *1 134.5,73 PMOS
M$45 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $46 r0 *1 137.5,73 PMOS
M$46 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $47 r0 *1 140.5,73 PMOS
M$47 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $48 r0 *1 143.5,73 PMOS
M$48 1 2 3 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $49 r0 *1 146.5,73 PMOS
M$49 3 2 1 4 PMOS L=1U W=140U AS=140P AD=140P PS=142U PD=142U
* device instance $50 r0 *1 149.5,73 PMOS
M$50 1 2 3 4 PMOS L=1U W=140U AS=140P AD=280P PS=142U PD=284U
.ENDS Pch$6

* cell Pch$7
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch$7 1 2 3 4
* device instance $1 r0 *1 2.5,23 PMOS
M$1 3 2 1 4 PMOS L=1U W=40U AS=80P AD=40P PS=84U PD=42U
* device instance $2 r0 *1 5.5,23 PMOS
M$2 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $3 r0 *1 8.5,23 PMOS
M$3 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $4 r0 *1 11.5,23 PMOS
M$4 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $5 r0 *1 14.5,23 PMOS
M$5 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $6 r0 *1 17.5,23 PMOS
M$6 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $7 r0 *1 20.5,23 PMOS
M$7 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $8 r0 *1 23.5,23 PMOS
M$8 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $9 r0 *1 26.5,23 PMOS
M$9 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $10 r0 *1 29.5,23 PMOS
M$10 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $11 r0 *1 32.5,23 PMOS
M$11 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $12 r0 *1 35.5,23 PMOS
M$12 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $13 r0 *1 38.5,23 PMOS
M$13 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $14 r0 *1 41.5,23 PMOS
M$14 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $15 r0 *1 44.5,23 PMOS
M$15 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $16 r0 *1 47.5,23 PMOS
M$16 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $17 r0 *1 50.5,23 PMOS
M$17 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $18 r0 *1 53.5,23 PMOS
M$18 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $19 r0 *1 56.5,23 PMOS
M$19 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $20 r0 *1 59.5,23 PMOS
M$20 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $21 r0 *1 62.5,23 PMOS
M$21 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $22 r0 *1 65.5,23 PMOS
M$22 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $23 r0 *1 68.5,23 PMOS
M$23 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $24 r0 *1 71.5,23 PMOS
M$24 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $25 r0 *1 74.5,23 PMOS
M$25 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $26 r0 *1 77.5,23 PMOS
M$26 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $27 r0 *1 80.5,23 PMOS
M$27 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $28 r0 *1 83.5,23 PMOS
M$28 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $29 r0 *1 86.5,23 PMOS
M$29 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $30 r0 *1 89.5,23 PMOS
M$30 1 2 3 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $31 r0 *1 92.5,23 PMOS
M$31 3 2 1 4 PMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $32 r0 *1 95.5,23 PMOS
M$32 1 2 3 4 PMOS L=1U W=40U AS=40P AD=80P PS=42U PD=84U
.ENDS Pch$7

* cell Nch$6
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$6 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 2.5,23 NMOS
M$1 1 3 2 4 NMOS L=1U W=40U AS=80P AD=40P PS=84U PD=42U
* device instance $2 r0 *1 5.5,23 NMOS
M$2 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $3 r0 *1 8.5,23 NMOS
M$3 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $4 r0 *1 11.5,23 NMOS
M$4 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $5 r0 *1 14.5,23 NMOS
M$5 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $6 r0 *1 17.5,23 NMOS
M$6 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $7 r0 *1 20.5,23 NMOS
M$7 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $8 r0 *1 23.5,23 NMOS
M$8 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $9 r0 *1 26.5,23 NMOS
M$9 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $10 r0 *1 29.5,23 NMOS
M$10 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $11 r0 *1 32.5,23 NMOS
M$11 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $12 r0 *1 35.5,23 NMOS
M$12 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $13 r0 *1 38.5,23 NMOS
M$13 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $14 r0 *1 41.5,23 NMOS
M$14 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $15 r0 *1 44.5,23 NMOS
M$15 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $16 r0 *1 47.5,23 NMOS
M$16 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $17 r0 *1 50.5,23 NMOS
M$17 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $18 r0 *1 53.5,23 NMOS
M$18 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $19 r0 *1 56.5,23 NMOS
M$19 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $20 r0 *1 59.5,23 NMOS
M$20 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $21 r0 *1 62.5,23 NMOS
M$21 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $22 r0 *1 65.5,23 NMOS
M$22 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $23 r0 *1 68.5,23 NMOS
M$23 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $24 r0 *1 71.5,23 NMOS
M$24 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $25 r0 *1 74.5,23 NMOS
M$25 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $26 r0 *1 77.5,23 NMOS
M$26 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $27 r0 *1 80.5,23 NMOS
M$27 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $28 r0 *1 83.5,23 NMOS
M$28 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $29 r0 *1 86.5,23 NMOS
M$29 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $30 r0 *1 89.5,23 NMOS
M$30 2 3 1 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $31 r0 *1 92.5,23 NMOS
M$31 1 3 2 4 NMOS L=1U W=40U AS=40P AD=40P PS=42U PD=42U
* device instance $32 r0 *1 95.5,23 NMOS
M$32 2 3 1 4 NMOS L=1U W=40U AS=40P AD=80P PS=42U PD=84U
.ENDS Nch$6
