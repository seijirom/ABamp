* Created by KLayout

* cell amp_ab
* pin VSS_P
* pin VDD_P
* pin TSD_IN
* pin SIGNAL_IN
* pin VDD
* pin CAP_G
* pin GND
.SUBCKT amp_ab 1 2 6 9 10 22 31
* net 1 VSS_P
* net 2 VDD_P
* net 6 TSD_IN
* net 9 SIGNAL_IN
* net 10 VDD
* net 22 CAP_G
* net 31 GND
* device instance $1 r0 *1 20,2.5 HRES
R$1 6 10 120750 HRES
* device instance $2 m90 *1 215,-190 NMOS
M$2 1 12 3 31 NMOS L=1U W=8000U AS=8080P AD=8080P PS=8282U PD=8282U
* device instance $102 r0 *1 227,-208.5 PMOS
M$102 3 4 2 2 PMOS L=1U W=28000U AS=28280P AD=28280P PS=29694U PD=29694U
* device instance $802 r0 *1 146,15 PMOS
M$802 10 7 4 10 PMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $806 r0 *1 134,-32 NMOS
M$806 12 16 4 31 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $807 m90 *1 124,-32 NMOS
M$807 8 16 16 31 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $808 m90 *1 88.5,-33 CAP
C$808 11 4 1.248e-11 CAP
* device instance $809 m90 *1 148,-32 PMOS
M$809 4 13 12 4 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $810 r0 *1 165,-32 PMOS
M$810 17 13 13 17 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $811 r0 *1 -1.5,-33.5 HRES
R$811 10 9 23000 HRES
* device instance $812 r0 *1 9,-33.5 HRES
R$812 31 9 23000 HRES
* device instance $813 m90 *1 52,-44.5 NMOS
M$813 14 5 11 31 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $814 r180 *1 52,-23.5 NMOS
M$814 7 5 11 31 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $815 r0 *1 34,-44.5 NMOS
M$815 14 9 15 31 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $816 m0 *1 34,-23.5 NMOS
M$816 19 9 15 31 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $817 m0 *1 34,-79 NMOS
M$817 14 6 31 31 NMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $821 m0 *1 127,-79 NMOS
M$821 12 6 31 31 NMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $825 r180 *1 21,-79 NMOS
M$825 6 6 31 31 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $827 m0 *1 160.5,-79.5 NMOS
M$827 13 6 31 31 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $829 r180 *1 1,-79 NMOS
M$829 18 6 31 31 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $831 m90 *1 58.5,14.5 PMOS
M$831 10 19 7 10 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $833 r0 *1 -4,14.5 PMOS
M$833 10 18 18 10 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $835 r0 *1 122.5,15 PMOS
M$835 10 18 16 10 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $837 r0 *1 34.5,14.5 PMOS
M$837 10 19 19 10 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $839 m90 *1 191.5,89 HRES
R$839 3 5 126500 HRES
* device instance $840 m90 *1 139.5,119 HRES
R$840 22 5 11500 HRES
* device instance $851 r180 *1 78.5,85 PMOS
M$851 10 17 17 10 PMOS L=1U W=1280U AS=1320P AD=1320P PS=1386U PD=1386U
* device instance $883 m90 *1 77,138 NMOS
M$883 31 8 8 31 NMOS L=1U W=1280U AS=1320P AD=1320P PS=1386U PD=1386U
.ENDS amp_ab
