* Created by KLayout

* cell amp_ab
.SUBCKT amp_ab
* net 28 SUBSTRATE
* device instance $1 r0 *1 -1.11,-34.64 HRES
R$1 2 7 20000
* device instance $2 r0 *1 9.39,-34.64 HRES
R$2 28 7 20000
* device instance $3 r0 *1 20.39,2.86 HRES
R$3 5 2 120750
* device instance $9 r0 *1 141.91,117.55 HRES
R$9 29 3 10000
* device instance $15 r0 *1 191.91,147.55 HRES
R$15 1 3 110000
* device instance $16 m90 *1 215.39,-174.29 NMOS
M$16 28 10 1 28 NMOS L=1U W=8000U AS=8080P AD=8080P PS=8282U PD=8282U
* device instance $116 r0 *1 227.48,-208.59 PMOS
M$116 1 4 2 2 PMOS L=1U W=28000U AS=28280P AD=28280P PS=29694U PD=29694U
* device instance $816 r0 *1 146.39,15.36 PMOS
M$816 2 6 4 2 PMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $820 r0 *1 134.39,-31.64 NMOS
M$820 10 16 4 28 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $821 m90 *1 124.39,-31.64 NMOS
M$821 8 16 16 28 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $822 m90 *1 88.89,-32.14 CAP
C$822 9 4 1.04e-11
* device instance $823 m90 *1 148.39,-31.64 PMOS
M$823 4 11 10 4 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $824 r0 *1 164.39,-31.64 PMOS
M$824 17 11 11 17 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $825 m90 *1 52.39,-44.14 NMOS
M$825 12 3 9 28 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $826 r180 *1 52.39,-23.14 NMOS
M$826 6 3 9 28 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $827 r0 *1 34.39,-44.14 NMOS
M$827 12 7 13 28 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $828 m0 *1 34.39,-23.14 NMOS
M$828 15 7 13 28 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $829 m0 *1 34.39,-78.64 NMOS
M$829 12 5 28 28 NMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $833 m0 *1 127.39,-78.64 NMOS
M$833 10 5 28 28 NMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $837 r180 *1 21.39,-78.64 NMOS
M$837 5 5 28 28 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $839 m0 *1 160.89,-79.14 NMOS
M$839 11 5 28 28 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $841 r180 *1 1.39,-78.64 NMOS
M$841 14 5 28 28 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $843 r0 *1 -3.61,14.86 PMOS
M$843 2 14 14 2 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $845 m90 *1 58.89,14.86 PMOS
M$845 2 15 6 2 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $847 r0 *1 122.89,15.36 PMOS
M$847 2 14 16 2 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $849 r0 *1 34.89,14.86 PMOS
M$849 2 15 15 2 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $851 r180 *1 78.67,85.35 PMOS
M$851 2 17 17 2 PMOS L=1U W=1280U AS=1320P AD=1320P PS=1386U PD=1386U
* device instance $883 m90 *1 77.02,138.26 NMOS
M$883 28 8 8 28 NMOS L=1U W=1280U AS=1320P AD=1320P PS=1386U PD=1386U
.ENDS amp_ab
