* Z:\HOME\SEIJIROM\WORK\2021_9\ABAMP\HARUNA_AB_TB_.ASC
*V1 N001 0 3.3
*C1 N003 OUT 1000U
*V2 IN 0 SINE({VIN_DC+VOFF} 0.1 1K) AC 1 0
*C3 N002 0 100U
*RL N003 0 8
*V3 N002 0 {VIN_DC}
*XX1 N002 IN N001 OUT N001 0 HARUNA_AB_
*
* BLOCK SYMBOL DEFINITIONS
.SUBCKT HARUNA_AB_ CAP_G SIGNAL_IN VDD OUT VDD_P VSS_P
M24 N006 IN_ N010 0 NMOS L=4U W=8U
M23 N007 SIGNAL_IN N010 0 NMOS L=4U W=8U
M25 N010 N011 0 0 NMOS L=4U W=160U
M22 N003 N002 VDD VDD PMOS L=4U W=80U
M21 N002 N002 VDD VDD PMOS L=4U W=80U
M7 N005 N003 VDD VDD PMOS L=4U W=160U
M9 N013 N011 0 0 NMOS L=4U W=160U
M27 N011 N011 0 0 NMOS L=4U W=80U
M2 OUT N013 VSS_P 0 NMOS L=1U W=8000U
M3 N004 N004 VDD VDD PMOS L=1U W=1280U
M12 N012 N012 0 0 NMOS L=1U W=1280U
M11 N008 N008 N012 0 NMOS L=4U W=20U
M8 N005 N008 N013 0 NMOS L=4U W=20U
M6 N013 N009 N005 N005 PMOS L=4U W=20U
M4 N009 N009 N004 N004 PMOS L=4U W=20U
M1 OUT N005 VDD_P VDD_P PMOS L=1U W=28000U
M5 N009 N011 0 0 NMOS L=4U W=80U
M26 N001 N001 VDD VDD PMOS L=4U W=80U
M10 N008 N001 VDD VDD PMOS L=4U W=80U
R2 IN_ CAP_G 10K
R1 OUT IN_ 110K
R11 VDD SIGNAL_IN 20K
R12 SIGNAL_IN 0 20K
R22 VDD N011 117K
M13 N001 N011 0 0 NMOS L=4U W=80U
C1 N005 N006 12P
M14 N003 IN_ N006 0 NMOS L=4U W=8U
M15 N002 SIGNAL_IN N007 0 NMOS L=4U W=8U
.ENDS HARUNA_AB_

.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\SEIJIROM\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
.TRAN 30M
*.INCLUDE "./MODELS/OR1_MOS"
;AC DEC 100 1 100MEG
* .STEP PARAM CC 2P 8P 2P
.PARAM CC=6P
* .STEP PARAM NP 300 600 100?
.PARAM NP=100
.PARAM VIN_DC=1.65
* .STEP PARAM VOFF _0.1 0.1 0.025
.PARAM VOFF=0
.MEAS TRAN A MAX V(N003)
.BACKANNO
.GLOBAL 0
.END
