* Created by KLayout

* cell amp_ab
* pin VDD_P
* pin VSS_P
* pin OUT
* pin TSD_IN
* pin SIGNAL_IN
* pin VDD
* pin CAP_G
* pin GND
.SUBCKT amp_ab 1 2 3 5 9 10 21 31
* net 1 VDD_P
* net 2 VSS_P
* net 3 OUT
* net 5 TSD_IN
* net 9 SIGNAL_IN
* net 10 VDD
* net 21 CAP_G
* net 31 GND
* device instance $1 m90 *1 215,-174.5 NMOS
M$1 2 12 3 31 NMOS L=1U W=8000U AS=8080P AD=8080P PS=8282U PD=8282U
* device instance $101 r0 *1 227,-209 PMOS
M$101 3 6 1 1 PMOS L=1U W=28000U AS=28280P AD=28280P PS=29694U PD=29694U
* device instance $801 r0 *1 146,15 PMOS
M$801 10 7 6 10 PMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $805 r0 *1 134,-32 NMOS
M$805 12 17 6 31 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $806 m90 *1 124,-32 NMOS
M$806 8 17 17 31 NMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $807 m90 *1 88.5,-33 CAP
C$807 11 6 1.248e-11 CAP
* device instance $808 m90 *1 148,-32 PMOS
M$808 6 13 12 6 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $809 r0 *1 164,-32 PMOS
M$809 18 13 13 18 PMOS L=4U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $810 r0 *1 20,2.5 HRES
R$810 5 10 120750 HRES
* device instance $811 r0 *1 -1.5,-35 HRES
R$811 10 9 20000 HRES
* device instance $812 r0 *1 9,-35 HRES
R$812 31 9 20000 HRES
* device instance $813 m90 *1 52,-44.5 NMOS
M$813 14 4 11 31 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $814 r180 *1 52,-23.5 NMOS
M$814 7 4 11 31 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $815 r0 *1 34,-44.5 NMOS
M$815 14 9 19 31 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $816 m0 *1 34,-23.5 NMOS
M$816 16 9 19 31 NMOS L=4U W=8U AS=16P AD=16P PS=20U PD=20U
* device instance $817 m0 *1 34,-79 NMOS
M$817 14 5 31 31 NMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $821 m0 *1 127,-79 NMOS
M$821 12 5 31 31 NMOS L=4U W=160U AS=200P AD=200P PS=210U PD=210U
* device instance $825 r180 *1 21,-79 NMOS
M$825 5 5 31 31 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $827 m0 *1 160.5,-79.5 NMOS
M$827 13 5 31 31 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $829 r180 *1 1,-79 NMOS
M$829 15 5 31 31 NMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $831 m90 *1 58.5,14.5 PMOS
M$831 10 16 7 10 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $833 r0 *1 -4,14.5 PMOS
M$833 10 15 15 10 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $835 r0 *1 122.5,15 PMOS
M$835 10 15 17 10 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $837 r0 *1 34.5,14.5 PMOS
M$837 10 16 16 10 PMOS L=4U W=80U AS=120P AD=120P PS=126U PD=126U
* device instance $841 m90 *1 141.5,117.5 HRES
R$841 21 4 10000 HRES
* device instance $848 m90 *1 191.5,147.5 HRES
R$848 3 4 110000 HRES
* device instance $851 r180 *1 78.5,85 PMOS
M$851 10 18 18 10 PMOS L=1U W=1280U AS=1320P AD=1320P PS=1386U PD=1386U
* device instance $883 m90 *1 77,138 NMOS
M$883 31 8 8 31 NMOS L=1U W=1280U AS=1320P AD=1320P PS=1386U PD=1386U
.ENDS amp_ab
